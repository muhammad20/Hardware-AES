
module thirtytwobitxor(out, in1, in2);
input [32:0] in1;
input [32:0] in2;
output [32:0] out;

xor(out[0],in1[0],in2[0]);
xor(out[1],in1[1],in2[1]);
xor(out[2],in1[2],in2[2]);
xor(out[3],in1[3],in2[3]);
xor(out[4],in1[4],in2[4]);
xor(out[5],in1[5],in2[5]);
xor(out[6],in1[6],in2[6]);
xor(out[7],in1[7],in2[7]);
xor(out[8],in1[8],in2[8]);
xor(out[9],in1[9],in2[9]);
xor(out[10],in1[10],in2[10]);
xor(out[11],in1[11],in2[11]);
xor(out[12],in1[12],in2[12]);
xor(out[13],in1[13],in2[13]);
xor(out[14],in1[14],in2[14]);
xor(out[15],in1[15],in2[15]);
xor(out[16],in1[16],in2[16]);
xor(out[17],in1[17],in2[17]);
xor(out[18],in1[18],in2[18]);
xor(out[19],in1[19],in2[19]);
xor(out[20],in1[20],in2[20]);
xor(out[21],in1[21],in2[21]);
xor(out[22],in1[22],in2[22]);
xor(out[23],in1[23],in2[23]);
xor(out[24],in1[24],in2[24]);
xor(out[25],in1[25],in2[25]);
xor(out[26],in1[26],in2[26]);
xor(out[27],in1[27],in2[27]);
xor(out[28],in1[28],in2[28]);
xor(out[29],in1[29],in2[29]);
xor(out[30],in1[30],in2[30]);
xor(out[31],in1[31],in2[31]);
xor(out[32],in1[32],in2[32]);

endmodule
