
module AddRoundKey(prevState, nextState,w,round);
input  [127:0]prevState ;
input  [1919:0]w;
input [4:0]round;
output [127:0] nextState ;
wire [7:0] s [0:3][0:3];
wire [7:0] sNew[ 0:3][0:3];
wire [31:0] wo [0:59];
wire [31:0] temp0;
wire [31:0] temp1;
wire [31:0] temp2;
wire [31:0] temp3;
wire [31:0] sCol0;
wire [31:0] sCol1;
wire [31:0] sCol2;
wire [31:0] sCol3;
wire  [31:0] sNewCol0;
wire  [31:0] sNewCol1;
wire  [31:0] sNewCol2;
wire  [31:0] sNewCol3;

assign wo[59]=w[31:0];
assign wo[58]=w[63:32];
assign wo[57]=w[95:64];
assign wo[56]=w[127:96];
assign wo[55]=w[159:128];
assign wo[54]=w[191:160];
assign wo[53]=w[223:192];
assign wo[52]=w[255:224];
assign wo[51]=w[287:256];
assign wo[50]=w[319:288];
assign wo[49]=w[351:320];
assign wo[48]=w[383:352];
assign wo[47]=w[415:384];
assign wo[46]=w[447:416];
assign wo[45]=w[479:448];
assign wo[44]=w[511:480];
assign wo[43]=w[543:512];
assign wo[42]=w[575:544];
assign wo[41]=w[607:576];
assign wo[40]=w[639:608];
assign wo[39]=w[671:640];
assign wo[38]=w[703:672];
assign wo[37]=w[735:704];
assign wo[36]=w[767:736];
assign wo[35]=w[799:768];
assign wo[34]=w[831:800];
assign wo[33]=w[863:832];
assign wo[32]=w[895:864];
assign wo[31]=w[927:896];
assign wo[30]=w[959:928];
assign wo[29]=w[991:960];
assign wo[28]=w[1023:992];
assign wo[27]=w[1055:1024];
assign wo[26]=w[1087:1056];
assign wo[25]=w[1119:1088];
assign wo[24]=w[1151:1120];
assign wo[23]=w[1183:1152];
assign wo[22]=w[1215:1184];
assign wo[21]=w[1247:1216];
assign wo[20]=w[1279:1248];
assign wo[19]=w[1311:1280];
assign wo[18]=w[1343:1312];
assign wo[17]=w[1375:1344];
assign wo[16]=w[1407:1376];
assign wo[15]=w[1439:1408];
assign wo[14]=w[1471:1440];
assign wo[13]=w[1503:1472];
assign wo[12]=w[1535:1504];
assign wo[11]=w[1567:1536];
assign wo[10]=w[1599:1568];
assign wo[9]=w[1631:1600];
assign wo[8]=w[1663:1632];
assign wo[7]=w[1695:1664];
assign wo[6]=w[1727:1696];
assign wo[5]=w[1759:1728];
assign wo[4]=w[1791:1760];
assign wo[3]=w[1823:1792];
assign wo[2]=w[1855:1824];
assign wo[1]=w[1887:1856];
assign wo[0]=w[1919:1888];

assign s[3][3] = prevState[7:0];
assign s[3][2] = prevState[15:8];
assign s[3][1] = prevState[23:16];
assign s[3][0] = prevState[31:24];
assign s[2][3] = prevState[39:32];
assign s[2][2] = prevState[47:40];
assign s[2][1] = prevState[55:48];
assign s[2][0] = prevState[63:56];
assign s[1][3] = prevState[71:64];
assign s[1][2] = prevState[79:72];
assign s[1][1] = prevState[87:80];
assign s[1][0] = prevState[95:88];
assign s[0][3] = prevState[103:96];
assign s[0][2] = prevState[111:104];
assign s[0][1] = prevState[119:112];
assign s[0][0] = prevState[127:120];

assign  sCol3   [7:0] = s[3][3];
assign  sCol2   [7:0] = s[3][2];
assign  sCol1   [7:0] = s[3][1];
assign  sCol0   [7:0] = s[3][0];
assign  sCol3  [15:8] = s[2][3];
assign  sCol2  [15:8] = s[2][2];
assign  sCol1  [15:8] = s[2][1];
assign  sCol0  [15:8] = s[2][0];
assign  sCol3 [23:16] = s[1][3];
assign  sCol2 [23:16] = s[1][2];
assign  sCol1 [23:16] = s[1][1];
assign  sCol0 [23:16] = s[1][0];
assign  sCol3 [31:24] = s[0][3];
assign  sCol2 [31:24] = s[0][2];
assign  sCol1 [31:24] = s[0][1];
assign  sCol0 [31:24] = s[0][0];

assign temp0 = wo[4*round];
assign temp1 = wo[4*round+1];
assign temp2 = wo[4*round+2];
assign temp3 = wo[4*round+3];

thirtytwobitxor m1 (sNewCol0, temp0, sCol0);
thirtytwobitxor m2 (sNewCol1, temp1, sCol1);
thirtytwobitxor m3 (sNewCol2, temp2, sCol2);
thirtytwobitxor m4 (sNewCol3, temp3, sCol3);

assign  sNew[3][3] = sNewCol3   [7:0];
assign  sNew[3][2] = sNewCol2   [7:0];
assign  sNew[3][1] = sNewCol1   [7:0];
assign  sNew[3][0] = sNewCol0   [7:0];
assign  sNew[2][3] = sNewCol3  [15:8];
assign  sNew[2][2] = sNewCol2  [15:8];
assign  sNew[2][1] = sNewCol1  [15:8];
assign  sNew[2][0] = sNewCol0  [15:8];
assign  sNew[1][3] = sNewCol3 [23:16];
assign  sNew[1][2] = sNewCol2 [23:16];
assign  sNew[1][1] = sNewCol1 [23:16];
assign  sNew[1][0] = sNewCol0 [23:16];
assign  sNew[0][3] = sNewCol3 [31:24];
assign  sNew[0][2] = sNewCol2 [31:24];
assign  sNew[0][1] = sNewCol1 [31:24];
assign  sNew[0][0] = sNewCol0 [31:24];

assign  nextState[7:0] = sNew[3][3];
assign  nextState[15:8] = sNew[3][2];
assign  nextState[23:16] = sNew[3][1];
assign  nextState[31:24] = sNew[3][0];
assign  nextState[39:32] = sNew[2][3];
assign  nextState[47:40] = sNew[2][2];
assign  nextState[55:48] = sNew[2][1];
assign  nextState[63:56] = sNew[2][0];
assign  nextState[71:64] = sNew[1][3];
assign  nextState[79:72] = sNew[1][2];
assign  nextState[87:80] = sNew[1][1];
assign  nextState[95:88] = sNew[1][0];
assign  nextState[103:96] = sNew[0][3];
assign  nextState[111:104] = sNew[0][2];
assign  nextState[119:112] = sNew[0][1];
assign  nextState[127:120] = sNew[0][0];

endmodule